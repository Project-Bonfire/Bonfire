--Copyright (C) 2016 Siavoosh Payandeh Azad

library ieee;
use ieee.std_logic_1164.all;
--use IEEE.STD_LOGIC_ARITH.ALL;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity FIFO_credit_based is
    generic (
        DATA_WIDTH: integer := 32
    );
    port (  reset: in  std_logic;
            clk: in  std_logic;
            RX: in std_logic_vector(DATA_WIDTH-1 downto 0);

            valid_in: in std_logic;
            valid_in_vc: in std_logic;

            read_en_N : in std_logic;
            read_en_E : in std_logic;
            read_en_W : in std_logic;
            read_en_S : in std_logic;
            read_en_L : in std_logic;

            read_en_vc_N : in std_logic;
            read_en_vc_E : in std_logic;
            read_en_vc_W : in std_logic;
            read_en_vc_S : in std_logic;
            read_en_vc_L : in std_logic;

            credit_out: out std_logic;
            credit_out_vc: out std_logic;

            empty_out: out std_logic;
            empty_out_vc: out std_logic;

            Data_out: out std_logic_vector(DATA_WIDTH-1 downto 0);
            Data_out_vc: out std_logic_vector(DATA_WIDTH-1 downto 0)
    );
end FIFO_credit_based;

architecture behavior of FIFO_credit_based is
   signal read_pointer, read_pointer_in,  write_pointer, write_pointer_in: std_logic_vector(3 downto 0);
   signal full, empty: std_logic;
   signal read_en, write_en: std_logic;

   signal read_pointer_vc, read_pointer_in_vc,  write_pointer_vc, write_pointer_in_vc: std_logic_vector(3 downto 0);
   signal full_vc, empty_vc: std_logic;
   signal read_en_vc, write_en_vc: std_logic;

   signal FIFO_MEM_1, FIFO_MEM_1_in : std_logic_vector(DATA_WIDTH-1 downto 0);
   signal FIFO_MEM_2, FIFO_MEM_2_in : std_logic_vector(DATA_WIDTH-1 downto 0);
   signal FIFO_MEM_3, FIFO_MEM_3_in : std_logic_vector(DATA_WIDTH-1 downto 0);
   signal FIFO_MEM_4, FIFO_MEM_4_in : std_logic_vector(DATA_WIDTH-1 downto 0);

   signal FIFO_MEM_vc_1, FIFO_MEM_vc_1_in : std_logic_vector(DATA_WIDTH-1 downto 0);
   signal FIFO_MEM_vc_2, FIFO_MEM_vc_2_in : std_logic_vector(DATA_WIDTH-1 downto 0);
   signal FIFO_MEM_vc_3, FIFO_MEM_vc_3_in : std_logic_vector(DATA_WIDTH-1 downto 0);
   signal FIFO_MEM_vc_4, FIFO_MEM_vc_4_in : std_logic_vector(DATA_WIDTH-1 downto 0);


begin
 --------------------------------------------------------------------------------------------
--                           block diagram of the FIFO!


 --------------------------------------------------------------------------------------------
--  circular buffer structure
--                                   <--- WriteP
--              ---------------------------------
--              |   3   |   2   |   1   |   0   |
--              ---------------------------------
--                                   <--- readP
 --------------------------------------------------------------------------------------------

   process (clk, reset)begin
        if reset = '0' then
            read_pointer  <= "0001";
            write_pointer <= "0001";

            FIFO_MEM_1 <= (others=>'0');
            FIFO_MEM_2 <= (others=>'0');
            FIFO_MEM_3 <= (others=>'0');
            FIFO_MEM_4 <= (others=>'0');

            credit_out <= '0';

            read_pointer_vc  <= "0001";
            write_pointer_vc <= "0001";

            FIFO_MEM_vc_1 <= (others=>'0');
            FIFO_MEM_vc_2 <= (others=>'0');
            FIFO_MEM_vc_3 <= (others=>'0');
            FIFO_MEM_vc_4 <= (others=>'0');

            credit_out_vc <= '0';

        elsif clk'event and clk = '1' then
            write_pointer <= write_pointer_in;
            read_pointer  <=  read_pointer_in;
            credit_out <= '0';
            if write_en = '1' then
                --write into the memory
                  FIFO_MEM_1 <= FIFO_MEM_1_in;
                  FIFO_MEM_2 <= FIFO_MEM_2_in;
                  FIFO_MEM_3 <= FIFO_MEM_3_in;
                  FIFO_MEM_4 <= FIFO_MEM_4_in;
            end if;
            if read_en = '1' then
              credit_out <= '1';
            end if;


            write_pointer_vc <= write_pointer_in_vc;
            read_pointer_vc  <=  read_pointer_in_vc;
            credit_out_vc <= '0';
            if write_en_vc = '1' then
                --write into the memory
                  FIFO_MEM_vc_1 <= FIFO_MEM_vc_1_in;
                  FIFO_MEM_vc_2 <= FIFO_MEM_vc_2_in;
                  FIFO_MEM_vc_3 <= FIFO_MEM_vc_3_in;
                  FIFO_MEM_vc_4 <= FIFO_MEM_vc_4_in;
            end if;
            if read_en_vc = '1' then
              credit_out_vc <= '1';
            end if;
        end if;
    end process;

 -- anything below here is pure combinational

   -- combinatorial part
   process(RX, write_pointer, FIFO_MEM_1, FIFO_MEM_2, FIFO_MEM_3, FIFO_MEM_4)begin
      case( write_pointer ) is
          when "0001" => FIFO_MEM_1_in <= RX;         FIFO_MEM_2_in <= FIFO_MEM_2; FIFO_MEM_3_in <= FIFO_MEM_3; FIFO_MEM_4_in <= FIFO_MEM_4;
          when "0010" => FIFO_MEM_1_in <= FIFO_MEM_1; FIFO_MEM_2_in <= RX;         FIFO_MEM_3_in <= FIFO_MEM_3; FIFO_MEM_4_in <= FIFO_MEM_4;
          when "0100" => FIFO_MEM_1_in <= FIFO_MEM_1; FIFO_MEM_2_in <= FIFO_MEM_2; FIFO_MEM_3_in <= RX;         FIFO_MEM_4_in <= FIFO_MEM_4;
          when "1000" => FIFO_MEM_1_in <= FIFO_MEM_1; FIFO_MEM_2_in <= FIFO_MEM_2; FIFO_MEM_3_in <= FIFO_MEM_3; FIFO_MEM_4_in <= RX;
          when others => FIFO_MEM_1_in <= FIFO_MEM_1; FIFO_MEM_2_in <= FIFO_MEM_2; FIFO_MEM_3_in <= FIFO_MEM_3; FIFO_MEM_4_in <= FIFO_MEM_4;
      end case ;
   end process;

  process(read_pointer, FIFO_MEM_1, FIFO_MEM_2, FIFO_MEM_3, FIFO_MEM_4)begin
    case( read_pointer ) is
        when "0001" => Data_out <= FIFO_MEM_1;
        when "0010" => Data_out <= FIFO_MEM_2;
        when "0100" => Data_out <= FIFO_MEM_3;
        when "1000" => Data_out <= FIFO_MEM_4;
        when others => Data_out <= FIFO_MEM_1;
    end case ;
  end process;

  read_en <= (read_en_N or read_en_E or read_en_W or read_en_S or read_en_L) and not empty;
  empty_out <= empty;


  process(write_en, write_pointer)begin
    if write_en = '1'then
       write_pointer_in <= write_pointer(2 downto 0)&write_pointer(3);
    else
       write_pointer_in <= write_pointer;
    end if;
  end process;

  process(read_en, empty, read_pointer)begin
       if (read_en = '1' and empty = '0') then
           read_pointer_in <= read_pointer(2 downto 0)&read_pointer(3);
       else
           read_pointer_in <= read_pointer;
       end if;
  end process;

  process(full, valid_in) begin
     if valid_in = '1' and full ='0' then
         write_en <= '1';
     else
         write_en <= '0';
     end if;
  end process;

  process(write_pointer, read_pointer) begin
      if read_pointer = write_pointer  then
              empty <= '1';
      else
              empty <= '0';
      end if;
      --      if write_pointer = read_pointer>>1 then
      if write_pointer = read_pointer(0)&read_pointer(3 downto 1) then
              full <= '1';
      else
              full <= '0';
      end if;
  end process;


  -------------------------------------------------------------------------------
  ---           VC stuff
  ---
  -------------------------------------------------------------------------------

  process(RX, write_pointer_vc, FIFO_MEM_1, FIFO_MEM_2, FIFO_MEM_3, FIFO_MEM_4)begin
     case( write_pointer_vc ) is
         when "0001" => FIFO_MEM_vc_1_in <= RX;            FIFO_MEM_vc_2_in <= FIFO_MEM_vc_2; FIFO_MEM_vc_3_in <= FIFO_MEM_vc_3; FIFO_MEM_vc_4_in <= FIFO_MEM_vc_4;
         when "0010" => FIFO_MEM_vc_1_in <= FIFO_MEM_vc_1; FIFO_MEM_vc_2_in <= RX;            FIFO_MEM_vc_3_in <= FIFO_MEM_vc_3; FIFO_MEM_vc_4_in <= FIFO_MEM_vc_4;
         when "0100" => FIFO_MEM_vc_1_in <= FIFO_MEM_vc_1; FIFO_MEM_vc_2_in <= FIFO_MEM_vc_2; FIFO_MEM_vc_3_in <= RX;            FIFO_MEM_vc_4_in <= FIFO_MEM_vc_4;
         when "1000" => FIFO_MEM_vc_1_in <= FIFO_MEM_vc_1; FIFO_MEM_vc_2_in <= FIFO_MEM_vc_2; FIFO_MEM_vc_3_in <= FIFO_MEM_vc_3; FIFO_MEM_vc_4_in <= RX;
         when others => FIFO_MEM_vc_1_in <= FIFO_MEM_vc_1; FIFO_MEM_vc_2_in <= FIFO_MEM_vc_2; FIFO_MEM_vc_3_in <= FIFO_MEM_vc_3; FIFO_MEM_vc_4_in <= FIFO_MEM_vc_4;
     end case ;
  end process;

  process(read_pointer_vc, FIFO_MEM_vc_1, FIFO_MEM_vc_2, FIFO_MEM_vc_3, FIFO_MEM_vc_4)begin
   case( read_pointer_vc ) is
       when "0001" => Data_out_vc <= FIFO_MEM_vc_1;
       when "0010" => Data_out_vc <= FIFO_MEM_vc_2;
       when "0100" => Data_out_vc <= FIFO_MEM_vc_3;
       when "1000" => Data_out_vc <= FIFO_MEM_vc_4;
       when others => Data_out_vc <= FIFO_MEM_vc_1;
   end case ;
  end process;

  read_en_vc <= (read_en_vc_N or read_en_vc_E or read_en_vc_W or read_en_vc_S or read_en_vc_L) and not empty_vc;
  empty_out_vc <= empty_vc;


  process(write_en_vc, write_pointer_vc)begin
   if write_en_vc = '1'then
      write_pointer_in_vc <= write_pointer_vc(2 downto 0)&write_pointer_vc(3);
   else
      write_pointer_in_vc <= write_pointer_vc;
   end if;
  end process;

  process(read_en_vc, empty_vc, read_pointer_vc)begin
      if (read_en_vc = '1' and empty_vc = '0') then
          read_pointer_in_vc <= read_pointer_vc(2 downto 0)&read_pointer_vc(3);
      else
          read_pointer_in_vc <= read_pointer_vc;
      end if;
  end process;

  process(full_vc, valid_in_vc) begin
    if valid_in_vc = '1' and full_vc ='0' then
        write_en_vc <= '1';
    else
        write_en_vc <= '0';
    end if;
  end process;

  process(write_pointer_vc, read_pointer_vc) begin
     if read_pointer_vc = write_pointer_vc  then
             empty_vc <= '1';
     else
             empty_vc <= '0';
     end if;
     --      if write_pointer = read_pointer>>1 then
     if write_pointer_vc = read_pointer_vc(0)&read_pointer_vc(3 downto 1) then
             full_vc <= '1';
     else
             full_vc <= '0';
     end if;
  end process;


end;
